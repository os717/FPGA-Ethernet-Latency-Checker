`ifndef _NODE_DEF_H_
`define _NODE_DEF_H_

`define ETHERNET_TYPE_REQUEST {16'h1000}
`define ETHERNET_TYPE_REPLY   {16'h1001}

`endif